module example (
    ports
);
    
endmodule
always @() begin
    
end


//mkmkmkmkm
/*


*/


include "stdio.h"
include
